module cpusim();
logic clk, reset;

core cpu_sim(clk, reset);

initial begin


end
endmodule