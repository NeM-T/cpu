module rom(
input logic [31:0] rom_addr, 
output logic [31:0] rom_out);

logic [31:0]rom_data [32'hf:0];

initial begin
rom_data[0] <= 32'b0000000_00010_00001_000_00001_0110011; //add x1, x2, x1
rom_data[1] <= 32'b0000000_00010_00001_000_00001_0110011; //add x1, x2, x1
rom_data[2] <= 32'b0100000_00010_00001_000_00001_0110011; //sub x1, x2, x1
rom_data[3] <= 32'b0000000_00010_00001_110_00011_0110011; //or x1, x2, x3
rom_data[4] <= 32'b0000000_00010_00001_111_00011_0110011; //and x1, x2, x3
rom_data[5] <= 32'b0000000_00010_00001_010_00000_0100011; //sw x1
rom_data[6] <= 32'b0000000_00000_00001_010_00001_0000011; //lw x1
rom_data[7] <= 32'b0000000_00011_00001_000_00001_0010011; //addi x1, 3, x1
rom_data[8] <= 32'b0000000_00011_00001_000_00001_0010011; //addi x1, 3, x1
rom_data[9] <= 32'b0000000_00011_00001_000_00001_0010011; //addi x1, 3, x1
rom_data[10] <= 32'b0000000_00011_00001_000_00001_0010011; //addi x1, 3, x1
rom_data[11] <= 32'b0000000_00011_00001_000_00001_0010011; //addi x1, 3, x1
rom_data[12] <= 32'b0000000_00011_00001_000_00001_0010011; //addi x1, 3, x1
rom_data[13] <= 32'b0000000_00011_00001_000_00001_0010011; //addi x1, 3, x1
rom_data[14] <= 32'b0000000_00011_00001_000_00001_0010011; //addi x1, 3, x1
rom_data[15] <= 32'b0000000_00011_00001_000_00001_0010011; //addi x1, 3, x1
end

always_comb rom_out <= rom_data[rom_addr];
endmodule
